`timescale 1ns/10ps
module testbench_simple();
reg a,b,s;

